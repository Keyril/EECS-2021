module register (z, d, clk, enable);

input [31:0] z;
input [31:0] d;
input clk;
input enable;






endmodule
